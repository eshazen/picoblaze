---- non-zero words: 405
---- FILLING with 619 ----
--
-- Inferred program rom test for PicoBlaze
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity monitor is

  port (
    address     : in  std_logic_vector(11 downto 0);
    instruction : out std_logic_vector(17 downto 0);
    addr_2      : in  std_logic_vector(11 downto 0);
    wen         : in  std_logic;
    di          : in  std_logic_vector(17 downto 0);
    do          : out std_logic_vector(17 downto 0);
    clk         : in  std_logic);

end entity monitor;


architecture syn of monitor is
  -- N.B. (0 to nn) order needed otherwise data is backwards!
  type ram_type is array (0 to 1023 ) of std_logic_vector(19 downto 0);
  signal RAM : ram_type := (
    X"0108B",
    X"2D002",
    X"01002",
    X"2D004",
    X"20133",
    X"20118",
    X"0153E",
    X"20136",
    X"01801",
    X"2013B",
    X"1D508",
    X"32016",
    X"1D50D",
    X"3201B",
    X"1D520",
    X"3A009",
    X"1D81F",
    X"32009",
    X"20136",
    X"2E580",
    X"11801",
    X"22009",
    X"1D801",
    X"32009",
    X"19801",
    X"20136",
    X"22009",
    X"2017D",
    X"01000",
    X"2E080",
    X"2F800",
    X"01801",
    X"01900",
    X"01A21",
    X"0A080",
    X"1D000",
    X"32035",
    X"1D020",
    X"36029",
    X"11801",
    X"22022",
    X"11901",
    X"2E8A0",
    X"11A01",
    X"1D906",
    X"32035",
    X"0A080",
    X"1D000",
    X"32035",
    X"11801",
    X"1D020",
    X"3602E",
    X"22022",
    X"2F920",
    X"0B920",
    X"01A21",
    X"01B30",
    X"1D900",
    X"32066",
    X"0A8A0",
    X"06000",
    X"06110",
    X"06220",
    X"06330",
    X"0A580",
    X"11801",
    X"1D520",
    X"3205B",
    X"1D500",
    X"3205B",
    X"20147",
    X"3A049",
    X"22040",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"04050",
    X"22040",
    X"2E0B0",
    X"11B01",
    X"2E1B0",
    X"11B01",
    X"2E2B0",
    X"11B01",
    X"2E3B0",
    X"11B01",
    X"11A01",
    X"19901",
    X"22039",
    X"0B501",
    X"0355F",
    X"0B020",
    X"1D550",
    X"320EB",
    X"1D553",
    X"320DF",
    X"1D545",
    X"320D2",
    X"1D542",
    X"3208D",
    X"1D555",
    X"32084",
    X"1D557",
    X"3207F",
    X"1D54A",
    X"3207C",
    X"22006",
    X"01B01",
    X"01A2C",
    X"20176",
    X"22006",
    X"0B634",
    X"0B735",
    X"26760",
    X"200C9",
    X"36078",
    X"20183",
    X"2017D",
    X"22006",
    X"200AC",
    X"00480",
    X"20183",
    X"00470",
    X"20183",
    X"00460",
    X"20183",
    X"2017D",
    X"22006",
    X"2013B",
    X"00650",
    X"1D62B",
    X"3209D",
    X"1D63D",
    X"320A2",
    X"1D624",
    X"36078",
    X"200AC",
    X"36078",
    X"00470",
    X"20183",
    X"00460",
    X"20183",
    X"2017D",
    X"22006",
    X"200AC",
    X"36078",
    X"00A60",
    X"00B70",
    X"2208D",
    X"200AC",
    X"36078",
    X"2DA06",
    X"2DB08",
    X"2D60A",
    X"2D70C",
    X"2D80E",
    X"11A01",
    X"13B00",
    X"2208D",
    X"200C9",
    X"35000",
    X"00840",
    X"1480E",
    X"1480E",
    X"1480E",
    X"1480E",
    X"00740",
    X"14706",
    X"14706",
    X"14706",
    X"14706",
    X"200C9",
    X"35000",
    X"00540",
    X"1450E",
    X"1450E",
    X"04750",
    X"1440C",
    X"1440C",
    X"01600",
    X"04640",
    X"036C0",
    X"200C9",
    X"35000",
    X"04640",
    X"2013B",
    X"06000",
    X"25000",
    X"2013B",
    X"19520",
    X"39000",
    X"1D540",
    X"3D000",
    X"0353F",
    X"00450",
    X"06000",
    X"25000",
    X"1D003",
    X"36078",
    X"0B634",
    X"0B735",
    X"2D606",
    X"2D708",
    X"0B638",
    X"2D60A",
    X"0B639",
    X"2D60C",
    X"0B63A",
    X"2D60E",
    X"22006",
    X"01600",
    X"0183F",
    X"1D002",
    X"3A0E8",
    X"0B634",
    X"1D003",
    X"3A0E8",
    X"0B838",
    X"19801",
    X"2010A",
    X"2017D",
    X"22006",
    X"01600",
    X"01700",
    X"01810",
    X"1D002",
    X"3A0F5",
    X"0B634",
    X"0B735",
    X"1D003",
    X"3A0F5",
    X"0B838",
    X"200F7",
    X"22006",
    X"2D606",
    X"2D708",
    X"00470",
    X"20183",
    X"00460",
    X"20183",
    X"2017F",
    X"09405",
    X"20183",
    X"09404",
    X"20183",
    X"09403",
    X"20183",
    X"2017D",
    X"11601",
    X"13700",
    X"19801",
    X"3A006",
    X"220F7",
    X"00460",
    X"20183",
    X"2017F",
    X"2017F",
    X"0A460",
    X"20183",
    X"2017F",
    X"11601",
    X"19801",
    X"39000",
    X"0D60F",
    X"3610E",
    X"2017D",
    X"2210A",
    X"01B01",
    X"01A1E",
    X"20176",
    X"14580",
    X"20136",
    X"25000",
    X"2154D",
    X"2156F",
    X"2156E",
    X"21569",
    X"21574",
    X"2156F",
    X"21572",
    X"21520",
    X"21556",
    X"21531",
    X"2152E",
    X"21534",
    X"2150D",
    X"21500",
    X"21545",
    X"21572",
    X"21572",
    X"2156F",
    X"21572",
    X"2150D",
    X"21500",
    X"2B031",
    X"2B001",
    X"25000",
    X"09000",
    X"0D004",
    X"36136",
    X"2D501",
    X"25000",
    X"2013E",
    X"35000",
    X"2213B",
    X"011A7",
    X"09000",
    X"0D008",
    X"36145",
    X"19101",
    X"31000",
    X"2213F",
    X"09501",
    X"25000",
    X"19530",
    X"3A155",
    X"1D50A",
    X"3A158",
    X"19511",
    X"3A155",
    X"1150A",
    X"1D510",
    X"3A158",
    X"1952A",
    X"3A155",
    X"1150A",
    X"1D510",
    X"3A158",
    X"01500",
    X"1450E",
    X"25000",
    X"25000",
    X"2013B",
    X"20136",
    X"20147",
    X"39000",
    X"01507",
    X"20136",
    X"22159",
    X"00510",
    X"20147",
    X"3D000",
    X"00450",
    X"14406",
    X"14406",
    X"14406",
    X"14406",
    X"00500",
    X"20147",
    X"3D000",
    X"04450",
    X"25000",
    X"20159",
    X"00450",
    X"14406",
    X"14406",
    X"14406",
    X"14406",
    X"20159",
    X"04450",
    X"25000",
    X"24BA0",
    X"1D500",
    X"31000",
    X"20136",
    X"11A01",
    X"13B00",
    X"22176",
    X"0150D",
    X"22136",
    X"01520",
    X"22136",
    X"11530",
    X"22136",
    X"00540",
    X"1450E",
    X"1450E",
    X"1450E",
    X"1450E",
    X"2018F",
    X"20136",
    X"00540",
    X"0350F",
    X"2018F",
    X"20136",
    X"25000",
    X"1950A",
    X"3A192",
    X"11507",
    X"1153A",
    X"25000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000"
    );
begin

  process (clk) is
  begin  -- process
    if clk'event and clk = '1' then     -- rising clock edge
      instruction <= RAM(to_integer(unsigned(address)))(17 downto 0);
      if wen = '1' then
        RAM(to_integer(unsigned(addr_2))) <= B"00" & di;
      end if;
    end if;
  end process;

  do <= RAM(to_integer(unsigned(addr_2)))(17 downto 0);

end syn;
